module puerta_and(output wire y, input wire a, b, c); // Si es estructural output wire, si es behavioral output reg (instanciar un módulo)
  assign y = a & b & c;
endmodule